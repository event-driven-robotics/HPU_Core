-------------------------------------------------------------------------------
-- neuserial_core
-------------------------------------------------------------------------------

-- ------------------------------------------------------------------------------
-- 
--  Revision 1.1:  07/25/2018
--  - Added SpiNNlink capabilities
--    (M. Casti - IIT)
--    
-- ------------------------------------------------------------------------------

library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

library HPU_lib;
    use HPU_lib.aer_pkg.all;
    use HPU_lib.HPUComponents_pkg.all;

library neuserial_lib;
    use neuserial_lib.NSComponents_pkg.all;

library neuelab_lib;
    use neuelab_lib.NEComponents_pkg.all;

library datapath_lib;
    use datapath_lib.DPComponents_pkg.neuserial_PAER_arbiter;
	
library spinn_neu_if_lib;
	use spinn_neu_if_lib.spinn_neu_pkg.all;
	

--****************************
--   PORT DECLARATION
--****************************

entity neuserial_core is
    generic (
        -- -----------------------    
        -- PAER        
        C_RX_HAS_PAER             : boolean                       := true;
        C_RX_PAER_L_SENS_ID       : std_logic_vector(2 downto 0)  := "000";
        C_RX_PAER_R_SENS_ID       : std_logic_vector(2 downto 0)  := "000";
        C_RX_PAER_A_SENS_ID       : std_logic_vector(2 downto 0)  := "001";
        C_TX_HAS_PAER             : boolean                       := true;
        C_PAER_DSIZE              : natural range 1 to 29         := 24;
        -- -----------------------        
        -- HSSAER
        C_RX_HAS_HSSAER           : boolean                       := true;
        C_RX_HSSAER_N_CHAN        : natural range 1 to 4          := 3;
        C_RX_SAER0_L_SENS_ID      : std_logic_vector(2 downto 0)  := "000";
        C_RX_SAER1_L_SENS_ID      : std_logic_vector(2 downto 0)  := "000";
        C_RX_SAER2_L_SENS_ID      : std_logic_vector(2 downto 0)  := "000";
        C_RX_SAER3_L_SENS_ID      : std_logic_vector(2 downto 0)  := "000";        
        C_RX_SAER0_R_SENS_ID      : std_logic_vector(2 downto 0)  := "000";
        C_RX_SAER1_R_SENS_ID      : std_logic_vector(2 downto 0)  := "000";
        C_RX_SAER2_R_SENS_ID      : std_logic_vector(2 downto 0)  := "000";
        C_RX_SAER3_R_SENS_ID      : std_logic_vector(2 downto 0)  := "000";        
        C_RX_SAER0_A_SENS_ID      : std_logic_vector(2 downto 0)  := "001";
        C_RX_SAER1_A_SENS_ID      : std_logic_vector(2 downto 0)  := "001";
        C_RX_SAER2_A_SENS_ID      : std_logic_vector(2 downto 0)  := "001";
        C_RX_SAER3_A_SENS_ID      : std_logic_vector(2 downto 0)  := "001";
        C_TX_HAS_HSSAER           : boolean                       := true;
        C_TX_HSSAER_N_CHAN        : natural range 1 to 4          := 3;
        -- -----------------------        
        -- GTP
        C_RX_HAS_GTP              : boolean                       := true;
        C_GTP_RXUSRCLK2_PERIOD_NS : real                          := 6.4;        
        C_TX_HAS_GTP              : boolean                       := true;
        C_GTP_TXUSRCLK2_PERIOD_NS : real                          := 6.4;  
        C_GTP_DSIZE               : positive                      := 16;
        -- -----------------------                
        -- SPINNLINK
        C_RX_HAS_SPNNLNK          : boolean                       := true;
        C_TX_HAS_SPNNLNK          : boolean                       := true;
        C_PSPNNLNK_WIDTH      	  : natural range 1 to 32         := 32;
        -- -----------------------
        -- INTERCEPTION
        C_RX_LEFT_INTERCEPTION    : boolean                       := false;
        C_RX_RIGHT_INTERCEPTION   : boolean                       := false;
        C_RX_AUX_INTERCEPTION     : boolean                       := false;
        -- -----------------------
        -- SIMULATION
        C_SIM_TIME_COMPRESSION     : boolean                      := false   -- When "TRUE", simulation time is "compressed": frequencies of internal clock enables are speeded-up 
        
    );
    port (
        --
        -- Clocks & Reset
        ---------------------
        -- Resets
        nRst                      : in  std_logic;
        -- System Clock domain
        Clk_i                     : in  std_logic;
        Timing_i                  : in  time_tick;
        -- HSSAER Clocks domain
        Clk_hs_p                  : in  std_logic;
        Clk_hs_n                  : in  std_logic;
        Clk_ls_p                  : in  std_logic;
        Clk_ls_n                  : in  std_logic;
        
        --
        -- TX Interface
        ---------------------
        -- Parallel AER
        TxPaerAddr_o            : out std_logic_vector(C_PAER_DSIZE-1 downto 0);
        TxPaerReq_o             : out std_logic;
        TxPaerAck_i             : in  std_logic;
        -- HSSAER channels
        TxHssaer_o               : out std_logic_vector(0 to C_TX_HSSAER_N_CHAN-1);
        -- GTP lines

        --
        -- RX Left Interface
        ---------------------
        -- Parallel AER
        LRxPaerAddr_i           : in  std_logic_vector(C_PAER_DSIZE-1 downto 0);
        LRxPaerReq_i            : in  std_logic;
        LRxPaerAck_o            : out std_logic;
        -- HSSAER channels
        LRxHssaer_i              : in  std_logic_vector(0 to C_RX_HSSAER_N_CHAN-1);
        -- GTP lines
        LRxRxGtpAlignRequest_o   : out std_logic;
        LRxGtpRxUsrClk2_i        : in  std_logic;
        LRxSoftResetRx_o         : out  std_logic;                                          
        LRxGtpDataValid_o        : out std_logic;          
        LRxGtpRxuserrdy_o        : out std_logic;              
        LRxGtpRxdata_i           : in  std_logic_vector(C_GTP_DSIZE-1 downto 0);           
        LRxGtpRxchariscomma_i    : in  std_logic_vector((C_GTP_DSIZE/8)-1 downto 0);        
        LRxGtpRxcharisk_i        : in  std_logic_vector((C_GTP_DSIZE/8)-1 downto 0);        
        LRxGtpRxdisperr_i        : in  std_logic_vector((C_GTP_DSIZE/8)-1 downto 0);        
        LRxGtpRxnotintable_i     : in  std_logic_vector((C_GTP_DSIZE/8)-1 downto 0);            
        LRxGtpRxbyteisaligned_i  : in  std_logic;                                           
        LRxGtpRxbyterealign_i    : in  std_logic;         
        LRxGtpPllLock_i          : in  std_logic;                                           
        LRxGtpPllRefclklost_i    : in  std_logic;   
               
        --
        -- RX Right Interface
        ---------------------
        -- Parallel AER
        RRxPaerAddr_i             : in  std_logic_vector(C_PAER_DSIZE-1 downto 0);
        RRxPaerReq_i              : in  std_logic;
        RRxPaerAck_o              : out std_logic;
        -- HSSAER channels
        RRxHssaer_i              : in  std_logic_vector(0 to C_RX_HSSAER_N_CHAN-1);
        -- GTP lines
        RRxRxGtpAlignRequest_o   : out std_logic;
        RRxGtpRxUsrClk2_i        : in  std_logic;
        RRxSoftResetRx_o         : out  std_logic;                                          
        RRxGtpDataValid_o        : out std_logic;          
        RRxGtpRxuserrdy_o        : out std_logic;              
        RRxGtpRxdata_i           : in  std_logic_vector(C_GTP_DSIZE-1 downto 0);           
        RRxGtpRxchariscomma_i    : in  std_logic_vector((C_GTP_DSIZE/8)-1 downto 0);        
        RRxGtpRxcharisk_i        : in  std_logic_vector((C_GTP_DSIZE/8)-1 downto 0);        
        RRxGtpRxdisperr_i        : in  std_logic_vector((C_GTP_DSIZE/8)-1 downto 0);        
        RRxGtpRxnotintable_i     : in  std_logic_vector((C_GTP_DSIZE/8)-1 downto 0);            
        RRxGtpRxbyteisaligned_i  : in  std_logic;                                           
        RRxGtpRxbyterealign_i    : in  std_logic;         
        RRxGtpPllLock_i          : in  std_logic;                                           
        RRxGtpPllRefclklost_i    : in  std_logic;   
               
        --
        -- Aux Interface
        ---------------------
        -- Parallel AER
        AuxRxPaerAddr_i           : in  std_logic_vector(C_PAER_DSIZE-1 downto 0);
        AuxRxPaerReq_i            : in  std_logic;
        AuxRxPaerAck_o            : out std_logic;
        -- HSSAER channels 
        AuxRxHssaer_i              : in  std_logic_vector(C_RX_HSSAER_N_CHAN-1 downto 0);
        -- GTP lines
        AuxRxRxGtpAlignRequest_o   : out std_logic;
        AuxRxGtpRxUsrClk2_i        : in  std_logic;
        AuxRxSoftResetRx_o         : out  std_logic;                                          
        AuxRxGtpDataValid_o        : out std_logic;          
        AuxRxGtpRxuserrdy_o        : out std_logic;              
        AuxRxGtpRxdata_i           : in  std_logic_vector(C_GTP_DSIZE-1 downto 0);           
        AuxRxGtpRxchariscomma_i    : in  std_logic_vector((C_GTP_DSIZE/8)-1 downto 0);        
        AuxRxGtpRxcharisk_i        : in  std_logic_vector((C_GTP_DSIZE/8)-1 downto 0);        
        AuxRxGtpRxdisperr_i        : in  std_logic_vector((C_GTP_DSIZE/8)-1 downto 0);        
        AuxRxGtpRxnotintable_i     : in  std_logic_vector((C_GTP_DSIZE/8)-1 downto 0);            
        AuxRxGtpRxbyteisaligned_i  : in  std_logic;                                           
        AuxRxGtpRxbyterealign_i    : in  std_logic;         
        AuxRxGtpPllLock_i          : in  std_logic;                                           
        AuxRxGtpPllRefclklost_i    : in  std_logic;   
               
        --
        -- SpiNNlink Interface
        ---------------------
        -- input SpiNNaker link interface
        LRxData2of7FromSpinnaker_i       : in  std_logic_vector(6 downto 0); 
        LRxAckToSpinnaker_o              : out std_logic;
        RRxData2of7FromSpinnaker_i       : in  std_logic_vector(6 downto 0); 
        RRxAckToSpinnaker_o              : out std_logic;
        AuxRxData2of7FromSpinnaker_i     : in  std_logic_vector(6 downto 0); 
        AuxRxAckToSpinnaker_o            : out std_logic;
        -- output SpiNNaker link interface
        TxData2of7ToSpinnaker_o          : out std_logic_vector(6 downto 0);
        TxAckFromSpinnaker_i             : in  std_logic;

        --
        -- FIFOs interfaces
        ---------------------
        FifoCoreDat_o             : out std_logic_vector(31 downto 0);
        FifoCoreRead_i            : in  std_logic;
        FifoCoreEmpty_o           : out std_logic;
        FifoCoreAlmostEmpty_o     : out std_logic;
        FifoCoreBurstReady_o      : out std_logic;
        FifoCoreFull_o            : out std_logic;
        FifoCoreNumData_o         : out std_logic_vector(10 downto 0);

        --
        CoreFifoDat_i             : in  std_logic_vector(31 downto 0);
        CoreFifoWrite_i           : in  std_logic;
        CoreFifoFull_o            : out std_logic;
        CoreFifoAlmostFull_o      : out std_logic;
        CoreFifoEmpty_o           : out std_logic;

        -----------------------------------------------------------------------
        -- uController Interface
        ---------------------
        -- Control
        CleanTimer_i              : in  std_logic;
        FlushRXFifos_i            : in  std_logic;
        FlushTXFifos_i            : in  std_logic;        
        --TxEnable_i              : in  std_logic;
        --TxPaerFlushFifos_i      : in  std_logic;
        --LRxEnable_i             : in  std_logic;
        --RRxEnable_i             : in  std_logic;
        LRxPaerFlushFifos_i       : in  std_logic;
        RRxPaerFlushFifos_i       : in  std_logic;
        AuxRxPaerFlushFifos_i     : in  std_logic;
        FullTimestamp_i           : in  std_logic;

        -- Configurations
        DmaLength_i               : in  std_logic_vector(15 downto 0);
        RemoteLoopback_i          : in  std_logic;
        LocNearLoopback_i         : in  std_logic;
        LocFarLPaerLoopback_i     : in  std_logic;
        LocFarRPaerLoopback_i     : in  std_logic;
        LocFarAuxPaerLoopback_i   : in  std_logic;
        LocFarLSaerLoopback_i     : in  std_logic;
        LocFarRSaerLoopback_i     : in  std_logic;
        LocFarAuxSaerLoopback_i   : in  std_logic;
        LocFarSaerLpbkCfg_i       : in  t_XConCfg;
        LocFarSpnnLnkLoopbackSel_i : in  std_logic_vector(1 downto 0);

        TxPaerEn_i                : in  std_logic;
        TxHSSaerEn_i              : in  std_logic;
        TxGtpEn_i                 : in  std_logic;
        TxSpnnLnkEn_i             : in  std_logic;
        TxDestSwitch_i            : in  std_logic_vector(2 downto 0);
        --TxPaerIgnoreFifoFull_i  : in  std_logic;
        TxPaerReqActLevel_i       : in  std_logic;
        TxPaerAckActLevel_i       : in  std_logic;
        TxSaerChanEn_i            : in  std_logic_vector(C_TX_HSSAER_N_CHAN-1 downto 0);
        --TxSaerChanCfg_i         : in  t_hssaerCfg_array(C_TX_HSSAER_N_CHAN-1 downto 0);

        -- TX Timestamp
        TxTSMode_i                : in  std_logic_vector(1 downto 0);
        TxTSTimeoutSel_i          : in  std_logic_vector(3 downto 0);
        TxTSRetrigCmd_i           : in  std_logic;
        TxTSRearmCmd_i            : in  std_logic;
        TxTSRetrigStatus_o        : out std_logic;
        TxTSTimeoutCounts_o       : out std_logic;
        TxTSMaskSel_i             : in  std_logic_vector(1 downto 0);
        
        --
        LRxPaerEn_i               : in  std_logic;
        RRxPaerEn_i               : in  std_logic;
        AuxRxPaerEn_i             : in  std_logic;
        LRxHSSaerEn_i             : in  std_logic;
        RRxHSSaerEn_i             : in  std_logic;
        AuxRxHSSaerEn_i           : in  std_logic;
        LRxGtpEn_i                : in  std_logic;
        RRxGtpEn_i                : in  std_logic;
        AuxRxGtpEn_i              : in  std_logic;
        LRxSpnnLnkEn_i            : in  std_logic;
        RRxSpnnLnkEn_i            : in  std_logic;
        AuxRxSpnnLnkEn_i          : in  std_logic;
        LRxSaerChanEn_i           : in  std_logic_vector(C_RX_HSSAER_N_CHAN-1 downto 0);
        RRxSaerChanEn_i           : in  std_logic_vector(C_RX_HSSAER_N_CHAN-1 downto 0);
        AuxRxSaerChanEn_i         : in  std_logic_vector(C_RX_HSSAER_N_CHAN-1 downto 0);
        RxPaerReqActLevel_i       : in  std_logic;
        RxPaerAckActLevel_i       : in  std_logic;
        RxPaerIgnoreFifoFull_i    : in  std_logic;
        RxPaerAckSetDelay_i       : in  std_logic_vector(7 downto 0);
        RxPaerSampleDelay_i       : in  std_logic_vector(7 downto 0);
        RxPaerAckRelDelay_i       : in  std_logic_vector(7 downto 0);

        -- Status
        WrapDetected_o            : out   std_logic;

        --TxPaerFifoEmpty_o       : out std_logic;
        TxSaerStat_o              : out t_TxSaerStat_array(C_TX_HSSAER_N_CHAN-1 downto 0);

		    LRxPaerFifoFull_o         : out std_logic;
		    RRxPaerFifoFull_o         : out std_logic;
		    AuxRxPaerFifoFull_o       : out std_logic;
        LRxSaerStat_o             : out t_RxSaerStat_array(C_RX_HSSAER_N_CHAN-1 downto 0);
        RRxSaerStat_o             : out t_RxSaerStat_array(C_RX_HSSAER_N_CHAN-1 downto 0);
        AUXRxSaerStat_o           : out t_RxSaerStat_array(C_RX_HSSAER_N_CHAN-1 downto 0);
        LRxGtpStat_o              : out t_RxGtpStat;
        RRxGtpStat_o              : out t_RxGtpStat;
        AUXRxGtpStat_o            : out t_RxGtpStat;
        TxSpnnlnkStat_o           : out t_TxSpnnlnkStat;
        LRxSpnnlnkStat_o          : out t_RxSpnnlnkStat;
        RRxSpnnlnkStat_o          : out t_RxSpnnlnkStat;
        AuxRxSpnnlnkStat_o        : out t_RxSpnnlnkStat;
    
        Spnn_start_key_i          : in  std_logic_vector(31 downto 0);  -- SpiNNaker "START to send data" command key
        Spnn_stop_key_i           : in  std_logic_vector(31 downto 0);  -- SpiNNaker "STOP to send data" command key
        Spnn_tx_mask_i            : in  std_logic_vector(31 downto 0);  -- SpiNNaker TX Data Mask
        Spnn_rx_mask_i            : in  std_logic_vector(31 downto 0);  -- SpiNNaker RX Data Mask 
        Spnn_ctrl_i               : in  std_logic_vector(31 downto 0);  -- SpiNNaker Control register 
        Spnn_status_o             : out std_logic_vector(31 downto 0);  -- SpiNNaker Status Register  

        --
        -- INTERCEPTION
        ---------------------
        RRxData_o                 : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        RRxSrcRdy_o               : out std_logic;
        RRxDstRdy_i               : in  std_logic;
        RRxBypassData_i           : in  std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        RRxBypassSrcRdy_i         : in  std_logic;
        RRxBypassDstRdy_o         : out std_logic;
        --
        LRxData_o                 : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        LRxSrcRdy_o               : out std_logic;
        LRxDstRdy_i               : in  std_logic;
        LRxBypassData_i           : in  std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        LRxBypassSrcRdy_i         : in  std_logic;
        LRxBypassDstRdy_o         : out std_logic;
        --
        AuxRxData_o               : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        AuxRxSrcRdy_o             : out std_logic;
        AuxRxDstRdy_i             : in  std_logic;
        AuxRxBypassData_i         : in  std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        AuxRxBypassSrcRdy_i       : in  std_logic;
        AuxRxBypassDstRdy_o       : out std_logic;        
        
        --
        -- LED drivers
        ---------------------
        LEDo_o                    : out std_logic;
        LEDr_o                    : out std_logic;
        LEDy_o                    : out std_logic;

        --
        -- DEBUG SIGNALS
        ---------------------
        DBG_dataOk                : out std_logic;

        DBG_din                   : out std_logic_vector(63 downto 0);     
        DBG_wr_en                 : out std_logic;  
        DBG_rd_en                 : out std_logic;     
        DBG_dout                  : out std_logic_vector(63 downto 0);          
        DBG_full                  : out std_logic;    
        DBG_almost_full           : out std_logic;    
        DBG_overflow              : out std_logic;       
        DBG_empty                 : out std_logic;           
        DBG_almost_empty          : out std_logic;    
        DBG_underflow             : out std_logic;     
        DBG_data_count            : out std_logic_vector(10 downto 0);
        DBG_CH0_DATA              : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        DBG_CH0_SRDY              : out std_logic;   
        DBG_CH0_DRDY              : out std_logic;        
        DBG_CH1_DATA              : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        DBG_CH1_SRDY              : out std_logic;   
        DBG_CH1_DRDY              : out std_logic;        
        DBG_CH2_DATA              : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        DBG_CH2_SRDY              : out std_logic;   
        DBG_CH2_DRDY              : out std_logic;
        DBG_Timestamp_xD          : out std_logic_vector(31 downto 0);
        DBG_MonInAddr_xD          : out std_logic_vector(31 downto 0);
        DBG_MonInSrcRdy_xS        : out std_logic;
        DBG_MonInDstRdy_xS        : out std_logic;
        DBG_RESETFIFO             : out std_logic;
        DBG_src_rdy               : out std_logic_vector(C_RX_HSSAER_N_CHAN-1 downto 0);
        DBG_dst_rdy               : out std_logic_vector(C_RX_HSSAER_N_CHAN-1 downto 0);
        DBG_err                   : out std_logic_vector(C_RX_HSSAER_N_CHAN-1 downto 0);  
        DBG_run                   : out std_logic_vector(C_RX_HSSAER_N_CHAN-1 downto 0);
        DBG_RX                    : out std_logic_vector(C_RX_HSSAER_N_CHAN-1 downto 0);
        DBG_FIFO_0                : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        DBG_FIFO_1                : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        DBG_FIFO_2                : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        DBG_FIFO_3                : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
        DBG_FIFO_4                : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0)
    );
-- translate_off
begin
    -- check the consistency of the generics
    assert (C_INTERNAL_DSIZE >= (C_PAER_DSIZE+3))
        report  "C_PAER_DSIZE should be at least " & string(integer'image(C_INTERNAL_DSIZE-4)) & "with current value" & CR &
                "of C_INTERNAL_DSIZE constant (see package aer_pkg)"
        severity failure;
-- translate_on
end entity neuserial_core;


--****************************
--   IMPLEMENTATION
--****************************

architecture str of neuserial_core is

    -----------------------------------------------------------------------------
    -- constants
    -----------------------------------------------------------------------------
    --
    -- this is the number of cycles the level on req has to be stable in order for
    -- a value change to be detected (and not interpreted as a possible glitch)
    --constant c_ReqStableCycles                      : positive := 31;
    --
    --constant c_SIFReqDelayCycles                    : natural  := 2;
    --constant c_SIFAckStableCycles                   : natural  := 3;
    --
    --constant c_DVS_SCX                              : boolean  := false;
    --
    constant c_TestEnableSequencerNoWait            : boolean  := false;
    constant c_TestEnableSequencerToMonitorLoopback : boolean  := false;
    constant c_EnableMonitorControlsSequencerToo    : boolean  := false;
    --
    --constant cTestEnableNoGaepButGenCounter        : boolean  := false;
    --constant c_LRxPaerHighBits : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  "0000";
    --constant c_LRxSaerHighBits : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  "0100";
    --constant c_LRxGtpHighBits  : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  "1000";
    --constant c_RRxPaerHighBits : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  "0001";
    --constant c_RRxSaerHighBits : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  "0101";
    --constant c_RRxGtpHighBits  : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  "1001";

    constant c_RIGHT_EYE : std_logic_vector(1 downto 0) := "01";
    constant c_LEFT_EYE  : std_logic_vector(1 downto 0) := "00";
    constant c_AUX1      : std_logic_vector(1 downto 0) := "10";
    constant c_PAER_SRC  : std_logic_vector(1 downto 0) := "00";
    constant c_SAER_SRC  : std_logic_vector(1 downto 0) := "01";
    constant c_GTP_SRC   : std_logic_vector(1 downto 0) := "10";

    -- This header coding comes from AERsensorsMap.xlsx (svn version r12867)
    constant C_EVENT_TYPE_ADDRESS   : std_logic := '0';
    constant C_EVENT_TYPE_TIMESTAMP : std_logic := '1';
    constant C_RESERVED             : std_logic_vector(C_INTERNAL_DSIZE-C_PAER_DSIZE-4-1 downto 0) := (others => '0');
    constant C_SRC_ID_CAMERA        : std_logic_vector(2 downto 0) := "000";
    constant C_SRC_ID_AUX_SKIN_SENS : std_logic_vector(2 downto 0) := "001";
    constant C_SRC_ID_OTHER_SENS    : std_logic_vector(2 downto 0) := "X1X";
    constant c_zero_vect : std_logic_vector(C_INTERNAL_DSIZE-C_PAER_DSIZE-4-1 downto 0) := (others => '0');

    constant c_LRxPaerHighBits    : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_PAER_L_SENS_ID;
    constant c_LRxSaerHighBits0   : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_SAER0_L_SENS_ID;
    constant c_LRxSaerHighBits1   : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_SAER1_L_SENS_ID;
    constant c_LRxSaerHighBits2   : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_SAER2_L_SENS_ID;
    constant c_LRxSaerHighBits3   : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_SAER3_L_SENS_ID;
    constant c_LRxGtpHighBits     : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & "111";                
    constant c_RRxPaerHighBits    : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_PAER_R_SENS_ID; 
    constant c_RRxSaerHighBits0   : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_SAER0_R_SENS_ID;
    constant c_RRxSaerHighBits1   : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_SAER1_R_SENS_ID;
    constant c_RRxSaerHighBits2   : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_SAER2_R_SENS_ID;
    constant c_RRxSaerHighBits3   : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_SAER3_R_SENS_ID;
    constant c_RRxGtpHighBits     : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & "111";               
    constant c_AuxRxPaerHighBits  : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_PAER_A_SENS_ID; 
    constant c_AuxRxSaerHighBits0 : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_SAER0_A_SENS_ID;
    constant c_AuxRxSaerHighBits1 : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_SAER1_A_SENS_ID;
    constant c_AuxRxSaerHighBits2 : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_SAER2_A_SENS_ID;
    constant c_AuxRxSaerHighBits3 : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & C_RX_SAER3_A_SENS_ID;
    constant c_AuxRxGtpHighBits   : std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE) :=  C_EVENT_TYPE_ADDRESS & c_zero_vect & "111";               


    -----------------------------------------------------------------------------
    -- types
    -----------------------------------------------------------------------------


    -----------------------------------------------------------------------------
    -- signals
    -----------------------------------------------------------------------------
	signal	Rst				 : std_logic;
	
    signal  i_rxMonSrc       : t_PaerSrc_array(2 downto 0);
    signal  i_rxMonDst       : t_PaerDst_array(2 downto 0);

    signal  i_txSeqData      : std_logic_vector(31 downto 0);
    signal  i_txSeqSrcRdy    : std_logic;
    signal  i_txSeqDstRdy    : std_logic;

    signal  i_rxMonData      : std_logic_vector(31 downto 0);
    signal  i_rxMonSrcRdy    : std_logic;
    signal  i_rxMonDstRdy    : std_logic;

    signal  i_seqData        : std_logic_vector(31 downto 0);
    signal  i_seqSrcRdy      : std_logic;
    signal  i_seqDstRdy      : std_logic;

    signal  i_monData        : std_logic_vector(31 downto 0);
    signal  i_monSrcRdy      : std_logic;
    signal  i_monDstRdy      : std_logic;

    signal  i_TxPaerAddr   : std_logic_vector(C_PAER_DSIZE-1 downto 0);
    signal  i_TxPaerReq    : std_logic;
    signal  i_TxPaerAck    : std_logic;
    signal  ii_TxPaerReq   : std_logic;
    signal  ii_TxPaerAck   : std_logic;

    signal  i_LRxPaerAddr  : std_logic_vector(C_PAER_DSIZE-1 downto 0);
    signal  i_LRxPaerReq   : std_logic;
    signal  i_LRxPaerAck   : std_logic;
    signal  ii_LRxPaerReq  : std_logic;
    signal  ii_LRxPaerAck  : std_logic;

    signal  i_RRxPaerAddr  : std_logic_vector(C_PAER_DSIZE-1 downto 0);
    signal  i_RRxPaerReq   : std_logic;
    signal  i_RRxPaerAck   : std_logic;
    signal  ii_RRxPaerReq  : std_logic;
    signal  ii_RRxPaerAck  : std_logic;

    signal  i_AuxRxPaerAddr: std_logic_vector(C_PAER_DSIZE-1 downto 0);
    signal  i_AuxRxPaerReq : std_logic;
    signal  i_AuxRxPaerAck : std_logic;
    signal  ii_AuxRxPaerReq: std_logic;
    signal  ii_AuxRxPaerAck: std_logic;

    signal  i_TxHssaer      : std_logic_vector(0 to C_TX_HSSAER_N_CHAN-1);
    signal  i_LRxHssaer     : std_logic_vector(0 to C_RX_HSSAER_N_CHAN-1);
    signal  i_RRxHssaer     : std_logic_vector(0 to C_RX_HSSAER_N_CHAN-1);
    signal  i_AuxRxHssaer   : std_logic_vector(0 to C_RX_HSSAER_N_CHAN-1);
    
    signal  i_LRxData2of7FromSpinnaker          : std_logic_vector(6 downto 0);
    signal  i_LRxAckToSpinnaker                 : std_logic;
    signal  i_RRxData2of7FromSpinnaker          : std_logic_vector(6 downto 0);
    signal  i_RRxAckToSpinnaker                 : std_logic;
    signal  i_AuxRxData2of7FromSpinnaker        : std_logic_vector(6 downto 0);
    signal  i_AuxRxAckToSpinnaker               : std_logic;
    signal  i_TxData2of7ToSpinnaker            : std_logic_vector(6 downto 0);
    signal  i_TXAckFromSpinnaker               : std_logic;
    signal  i_Spnn_offload_on                   : std_logic;
    signal  i_Spnn_offload_off                  : std_logic;
    signal  i_Spnn_cmd_start                    : std_logic;
    signal  i_Spnn_cmd_stop                     : std_logic;

    signal  RRxData                             : std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
    signal  RRxSrcRdy                           : std_logic;
    signal  RRxDstRdy                           : std_logic;

    signal  LRxData                             : std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
    signal  LRxSrcRdy                           : std_logic;
    signal  LRxDstRdy                           : std_logic;

    signal  AuxRxData                           : std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
    signal  AuxRxSrcRdy                         : std_logic;
    signal  AuxRxDstRdy                         : std_logic;

--    for all : neuserial_loopback     use entity neuserial_lib.neuserial_loopback(beh);
--    for all : hpu_tx_datapath        use entity datapath_lib.hpu_tx_datapath(str);
--    for all : hpu_rx_datapath        use entity datapath_lib.hpu_rx_datapath(str);
--    for all : neuserial_PAER_arbiter use entity datapath_lib.neuserial_PAER_arbiter(rtl);
--    for all : CoreMonSeqRR           use entity neuelab_lib.CoreMonSeqRR(str);

-- GTP

-- --------------
-- GTP RX Left
signal i_LRxGtpRxDataRate     : std_logic_vector(15 downto 0);
signal i_LRxGtpRxAlignRate    : std_logic_vector( 7 downto 0);
signal i_LRxGtpRxMsgRate      : std_logic_vector(15 downto 0);
signal i_LRxGtpRxIdleRate     : std_logic_vector(15 downto 0);
signal i_LRxGtpRxEventRate    : std_logic_vector(15 downto 0);
signal i_LRxGtpRxMessageRate  : std_logic_vector( 7 downto 0);

-- GTP RX Right
signal i_RRxGtpRxDataRate     : std_logic_vector(15 downto 0);
signal i_RRxGtpRxAlignRate    : std_logic_vector( 7 downto 0);
signal i_RRxGtpRxMsgRate      : std_logic_vector(15 downto 0);
signal i_RRxGtpRxIdleRate     : std_logic_vector(15 downto 0);
signal i_RRxGtpRxEventRate    : std_logic_vector(15 downto 0);
signal i_RRxGtpRxMessageRate  : std_logic_vector( 7 downto 0);

-- GTP RX Aux
signal i_AuxRxGtpRxDataRate     : std_logic_vector(15 downto 0);
signal i_AuxRxGtpRxAlignRate    : std_logic_vector( 7 downto 0);
signal i_AuxRxGtpRxMsgRate      : std_logic_vector(15 downto 0);
signal i_AuxRxGtpRxIdleRate     : std_logic_vector(15 downto 0);
signal i_AuxRxGtpRxEventRate    : std_logic_vector(15 downto 0);
signal i_AuxRxGtpRxMessageRate  : std_logic_vector( 7 downto 0);

-- --------------
-- GTPTX




begin

	Rst <= not nRst;

    -- PAER Req and acknowledge polarity
    --
    TxPaerReq_o   <= ii_TxPaerReq  xnor TxPaerReqActLevel_i;
    ii_TxPaerAck  <= TxPaerAck_i   xnor TxPaerAckActLevel_i;

    ii_LRxPaerReq <= LRxPaerReq_i  xnor RxPaerReqActLevel_i;
    LRxPaerAck_o  <= ii_LRxPaerAck xnor RxPaerAckActLevel_i;

    ii_RRxPaerReq <= RRxPaerReq_i  xnor RxPaerReqActLevel_i;
    RRxPaerAck_o  <= ii_RRxPaerAck xnor RxPaerAckActLevel_i;

    ii_AuxRxPaerReq <= AuxRxPaerReq_i  xnor RxPaerReqActLevel_i;
    AuxRxPaerAck_o <= ii_AuxRxPaerAck xnor RxPaerAckActLevel_i;

    ------------------------
    -- Local Far Loopback
    ------------------------

    u_neuserial_loopback : neuserial_loopback
        generic map (
            C_PAER_DSIZE          => C_PAER_DSIZE,
            C_RX_HSSAER_N_CHAN    => C_RX_HSSAER_N_CHAN,
            C_TX_HSSAER_N_CHAN    => C_TX_HSSAER_N_CHAN
        )
        port map (
            Rx1PaerLpbkEn         => LocFarLPaerLoopback_i,      -- in  std_logic;
            Rx2PaerLpbkEn         => LocFarRPaerLoopback_i,      -- in  std_logic;
            Rx3PaerLpbkEn         => LocFarAuxPaerLoopback_i,    -- in  std_logic;
            Rx1SaerLpbkEn         => LocFarLSaerLoopback_i,      -- in  std_logic;
            Rx2SaerLpbkEn         => LocFarRSaerLoopback_i,      -- in  std_logic;
            Rx3SaerLpbkEn         => LocFarAuxSaerLoopback_i,    -- in  std_logic;
            XConSerCfg            => LocFarSaerLpbkCfg_i,        -- in  t_XConCfg;
            RxSpnnLnkLpbkEnSel    => LocFarSpnnLnkLoopbackSel_i, -- in  std_logic_vector(1 downto 0);

            -- Parallel AER
            ExtTxPAER_Addr_o      => TxPaerAddr_o,             -- out std_logic_vector(C_PAER_DSIZE-1 downto 0);
            ExtTxPAER_Req_o       => ii_TxPaerReq,             -- out std_logic;
            ExtTxPAER_Ack_i       => ii_TxPaerAck,             -- in  std_logic;

            ExtRx1PAER_Addr_i     => LRxPaerAddr_i,            -- in  std_logic_vector(C_PAER_DSIZE-1 downto 0);
            ExtRx1PAER_Req_i      => ii_LRxPaerReq,            -- in  std_logic;
            ExtRx1PAER_Ack_o      => ii_LRxPaerAck,            -- out std_logic;

            ExtRx2PAER_Addr_i     => RRxPaerAddr_i,            -- in  std_logic_vector(C_PAER_DSIZE-1 downto 0);
            ExtRx2PAER_Req_i      => ii_RRxPaerReq,            -- in  std_logic;
            ExtRx2PAER_Ack_o      => ii_RRxPaerAck,            -- out std_logic;

            ExtRx3PAER_Addr_i     => AuxRxPaerAddr_i,          -- in  std_logic_vector(C_PAER_DSIZE-1 downto 0);
            ExtRx3PAER_Req_i      => ii_AuxRxPaerReq,          -- in  std_logic;
            ExtRx3PAER_Ack_o      => ii_AuxRxPaerAck,          -- out std_logic;

            -- HSSAER
            ExtTxHSSAER_Tx_o      => TxHssaer_o,                -- out std_logic_vector(0 to C_TX_HSSAER_N_CHAN-1);
            ExtRx1HSSAER_Rx_i     => LRxHssaer_i,               -- in  std_logic_vector(0 to C_RX_HSSAER_N_CHAN-1);
            ExtRx2HSSAER_Rx_i     => RRxHssaer_i,               -- in  std_logic_vector(0 to C_RX_HSSAER_N_CHAN-1);
            ExtRx3HSSAER_Rx_i     => AuxRxHssaer_i,             -- in  std_logic_vector(0 to C_RX_HSSAER_N_CHAN-1);

            -- GTP interface
            --
            -- TBD signals to drive the GTP module
            --
            -- SpiNNlink interface
            ExtTx_data_2of7_to_spinnaker_o      => TxData2of7ToSpinnaker_o,     -- out std_logic_vector(6 downto 0);
            ExtTx_ack_from_spinnaker_i          => TxAckFromSpinnaker_i,         -- in  std_logic;
            ExtRx1_data_2of7_from_spinnaker_i   => LRxData2of7FromSpinnaker_i,  -- in  std_logic_vector(6 downto 0); 
            ExtRx1_ack_to_spinnaker_o           => LRxAckToSpinnaker_o,          -- out std_logic;
            ExtRx2_data_2of7_from_spinnaker_i   => RRxData2of7FromSpinnaker_i,  -- in  std_logic_vector(6 downto 0); 
            ExtRx2_ack_to_spinnaker_o           => RRxAckToSpinnaker_o,          -- out std_logic;
            ExtRx3_data_2of7_from_spinnaker_i   => AuxRxData2of7FromSpinnaker_i,-- in  std_logic_vector(6 downto 0); 
            ExtRx3_ack_to_spinnaker_o           => AuxRxAckToSpinnaker_o,        -- out std_logic;
            
          
            -- Parallel AER 
            CoreTxPAER_Addr_i     => i_TxPaerAddr,             -- in  std_logic_vector(C_PAER_DSIZE-1 downto 0);
            CoreTxPAER_Req_i      => i_TxPaerReq,              -- in  std_logic;
            CoreTxPAER_Ack_o      => i_TxPaerAck,              -- out std_logic;

            CoreRx1PAER_Addr_o    => i_LRxPaerAddr,            -- out std_logic_vector(C_PAER_DSIZE-1 downto 0);
            CoreRx1PAER_Req_o     => i_LRxPaerReq,             -- out std_logic;
            CoreRx1PAER_Ack_i     => i_LRxPaerAck,             -- in  std_logic;

            CoreRx2PAER_Addr_o    => i_RRxPaerAddr,            -- out std_logic_vector(C_PAER_DSIZE-1 downto 0);
            CoreRx2PAER_Req_o     => i_RRxPaerReq,             -- out std_logic;
            CoreRx2PAER_Ack_i     => i_RRxPaerAck,             -- in  std_logic;

            CoreRx3PAER_Addr_o    => i_AuxRxPaerAddr,          -- out std_logic_vector(C_PAER_DSIZE-1 downto 0);
            CoreRx3PAER_Req_o     => i_AuxRxPaerReq,           -- out std_logic;
            CoreRx3PAER_Ack_i     => i_AuxRxPaerAck,           -- in  std_logic;

            -- HSSAER
            CoreTxHSSAER_Tx_i     => i_TxHssaer,                -- in  std_logic_vector(0 to C_TX_HSSAER_N_CHAN-1);
            CoreRx1HSSAER_Rx_o    => i_LRxHssaer,               -- out std_logic_vector(0 to C_RX_HSSAER_N_CHAN-1);
            CoreRx2HSSAER_Rx_o    => i_RRxHssaer,               -- out std_logic_vector(0 to C_RX_HSSAER_N_CHAN-1);
            CoreRx3HSSAER_Rx_o    => i_AuxRxHssaer,             -- out std_logic_vector(0 to C_RX_HSSAER_N_CHAN-1)

            -- GTP interface
            --
            -- TBD signals to drive the GTP module
            --

            -- SpiNNlink interface
            CoreTx_data_2of7_to_spinnaker_i     => i_TxData2of7ToSpinnaker,     -- in  std_logic_vector(6 downto 0);
            CoreTx_ack_from_spinnaker_o         => i_TxAckFromSpinnaker,         -- out std_logic;
            CoreRx1_data_2of7_from_spinnaker_o  => i_LRxData2of7FromSpinnaker,  -- out std_logic_vector(6 downto 0); 
            CoreRx1_ack_to_spinnaker_i          => i_LRxAckToSpinnaker,          -- in  std_logic;
            CoreRx2_data_2of7_from_spinnaker_o  => i_RRxData2of7FromSpinnaker,  -- out std_logic_vector(6 downto 0); 
            CoreRx2_ack_to_spinnaker_i          => i_RRxAckToSpinnaker,          -- in  std_logic;
            CoreRx3_data_2of7_from_spinnaker_o  => i_AuxRxData2of7FromSpinnaker,-- out std_logic_vector(6 downto 0); 
            CoreRx3_ack_to_spinnaker_i          => i_AuxRxAckToSpinnaker         -- in  std_logic
        );

    
    ---------------------
    -- TX path
    ---------------------
    
    i_Spnn_offload_on  <= i_Spnn_cmd_stop or  Spnn_ctrl_i(2);
    i_Spnn_offload_off <= i_Spnn_cmd_start or Spnn_ctrl_i(1);

    u_tx_datapath : hpu_tx_datapath
        generic map (
            C_INPUT_DSIZE    => 32,
            C_PAER_DSIZE     => C_PAER_DSIZE,
            C_HAS_PAER       => C_TX_HAS_PAER,
            C_HAS_HSSAER     => C_TX_HAS_HSSAER,
            C_HSSAER_N_CHAN  => C_TX_HSSAER_N_CHAN,
            C_HAS_GTP        => C_TX_HAS_GTP,
            C_HAS_SPNNLNK    => C_TX_HAS_SPNNLNK,
            C_PSPNNLNK_WIDTH => C_PSPNNLNK_WIDTH
            
        )
        port map (
            -- Clocks & Reset
            nRst                 => nRst,                        -- in  std_logic;
            Clk_core             => Clk_i,                    -- in  std_logic;
			      Clk_ls_p             => Clk_ls_p,                     -- in  std_logic;
			      Clk_ls_n             => Clk_ls_n,                     -- in  std_logic;

            -----------------------------
            -- uController Interface
            -----------------------------

            -- Control signals
            -----------------------------
            --EnableIp_i           => TxEnable_i,                  -- in  std_logic;
			--PaerFlushFifos_i     => TxPaerFlushFifos_i,          -- in  std_logic;

            -- Status signals
            -----------------------------
            --PaerFifoFull_o       => TxPaerFifoEmpty_o,           -- out std_logic;
            TxSaerStat_o         => TxSaerStat_o,                -- out t_TxSaerStat_array(C_HSSAER_N_CHAN-1 downto 0);
            TxSpnnlnkStat_o      => TxSpnnlnkStat_o,             -- out t_TxSpnnlnkStat;
            
            -- Configuration signals
            -----------------------------
            --
            -- Destination I/F configurations
            EnablePAER_i         => TxPaerEn_i,                  -- in  std_logic;
            EnableHSSAER_i       => TxHSSaerEn_i,                -- in  std_logic;
            EnableGTP_i          => TxGtpEn_i,                   -- in  std_logic;
            EnableSPNNLNK_i      => TxSpnnLnkEn_i,
            DestinationSwitch_i  => TxDestSwitch_i,              -- in  std_logic_vector(2 downto 0);
            -- PAER
            --PaerIgnoreFifoFull_i => TxPaerIgnoreFifoFull_i,      -- in  std_logic;
            PaerReqActLevel_i    => '1',                         -- in  std_logic;
            PaerAckActLevel_i    => '1',                         -- in  std_logic;
            -- HSSAER
            HSSaerChanEn_i       => TxSaerChanEn_i,              -- in  std_logic_vector(C_HSSAER_N_CHAN-1 downto 0);
            --HSSAERChanCfg_i      => TxHSSaerChanCfg_i,           -- in  t_hssaerCfg_array(C_HSSAER_N_CHAN-1 downto 0);
            -- GTP
            --
            -- SpiNNaker
            -----------------------------
            Spnn_offload_on_i       => i_Spnn_offload_on,          -- in  std_logic;
            Spnn_offload_off_i      => i_Spnn_offload_off,         -- in  std_logic;            
            Spnn_tx_mask_i          => Spnn_tx_mask_i,             -- in  std_logic_vector(31 downto 0);
            Spnn_Offload_o          => Spnn_status_o(1),           -- out std_logic;
            Spnn_Link_Timeout_o     => Spnn_status_o(0),           -- out std_logic;
            Spnn_Link_Timeout_dis_i => Spnn_ctrl_i(0),             -- in  std_logic;       
                  
            -----------------------------
            -- Sequencer interface
            -----------------------------
            FromSeqDataIn_i      => i_txSeqData,                 -- in  std_logic_vector(C_INPUT_DSIZE-1 downto 0);
            FromSeqSrcRdy_i      => i_txSeqSrcRdy,               -- in  std_logic;
            FromSeqDstRdy_o      => i_txSeqDstRdy,               -- out std_logic;
        
            -----------------------------
            -- Destination interfaces
            -----------------------------
            -- Parallel AER
            PAER_Addr_o          => i_TxPaerAddr,              -- out std_logic_vector(C_PAER_DSIZE-1 downto 0);
            PAER_Req_o           => i_TxPaerReq,               -- out std_logic;
            PAER_Ack_i           => i_TxPaerAck,               -- in  std_logic;

            -- HSSAER
            HSSAER_Tx_o          => i_TxHssaer,                  -- out std_logic_vector(0 to C_HSSAER_N_CHAN-1)

            -- GTP interface
            --
            -- TBD signals to drive the GTP
            --

		    -- SpiNNlink 
		    data_2of7_to_spinnaker_o	=> i_TxData2of7ToSpinnaker,
		    ack_from_spinnaker_i      => i_TxAckFromSpinnaker

            -----------------------------
            -- Debug signals
            -----------------------------
        );
    
   
    
---------------------
-- RX paths
---------------------

u_rx_left_datapath : hpu_rx_datapath
  generic map (
    C_OUTPUT_DSIZE            => C_INTERNAL_DSIZE,
    C_PAER_DSIZE              => C_PAER_DSIZE,
    C_HAS_PAER                => C_RX_HAS_PAER,
    C_HAS_HSSAER              => C_RX_HAS_HSSAER,
    C_HSSAER_N_CHAN           => C_RX_HSSAER_N_CHAN,
    C_HAS_GTP                 => C_RX_HAS_GTP,
    C_GTP_DSIZE               => C_GTP_DSIZE,
    C_GTP_TXUSRCLK2_PERIOD_NS => C_GTP_TXUSRCLK2_PERIOD_NS,
    C_GTP_RXUSRCLK2_PERIOD_NS => C_GTP_RXUSRCLK2_PERIOD_NS,
    C_HAS_SPNNLNK             => C_RX_HAS_SPNNLNK,
    C_PSPNNLNK_WIDTH          => C_PSPNNLNK_WIDTH,
    C_SIM_TIME_COMPRESSION    => C_SIM_TIME_COMPRESSION
    )
  port map (

    -- **********************************************
    -- Barecontrol
    -- **********************************************
    -- Resets
    nRst                 => nRst,                         -- in  std_logic;
    -- System Clock domain
    Clk_i                => Clk_i,                        -- in  std_logic;
    En1Sec_i             => timing_i.en1s,                -- : in  std_logic;
		-- HSSAER Clocks domain
		Clk_hs_p             => Clk_hs_p,                     -- in  std_logic;
		Clk_hs_n             => Clk_hs_n,                     -- in  std_logic;
    Clk_ls_p             => Clk_ls_p,                     -- in  std_logic;
    Clk_ls_n             => Clk_ls_n,                     -- in  std_logic;
 
 
    -- **********************************************
    -- Controls
    -- **********************************************
    --
    -- In case of aux channel the HPU header is 
    -- adapted to what received
    -- ----------------------------------------------
    Aux_Channel_i        => '0',


    -- **********************************************
    -- uController Interface
    -- **********************************************

    -- Control signals
    -- ----------------------------------------------
    PaerFlushFifos_i     => LRxPaerFlushFifos_i,         -- in  std_logic;
    
    -- Status signals
    -----------------------------
    PaerFifoFull_o       => LRxPaerFifoFull_o,           -- out std_logic;
    RxSaerStat_o         => LRxSaerStat_o,               -- out t_RxSaerStat_array(C_HSSAER_N_CHAN-1 downto 0);
    RxGtpStat_o          => LRxGtpStat_o,                -- out t_RxGtpStat;
    RxSpnnlnkStat_o      => LRxSpnnlnkStat_o,            -- out t_RxSpnnlnkStat;
        
    -- GTP Statistics        
    GtpRxDataRate_o      => i_LRxGtpRxDataRate,           -- : out std_logic_vector(15 downto 0); -- Count per millisecond 
    GtpRxAlignRate_o     => i_LRxGtpRxAlignRate,          -- : out std_logic_vector( 7 downto 0); -- Count per millisecond 
    GtpRxMsgRate_o       => i_LRxGtpRxMsgRate,            -- : out std_logic_vector(15 downto 0); -- Count per millisecond 
    GtpRxIdleRate_o      => i_LRxGtpRxIdleRate,           -- : out std_logic_vector(15 downto 0); -- Count per millisecond 
    GtpRxEventRate_o     => i_LRxGtpRxEventRate,          -- : out std_logic_vector(15 downto 0); -- Count per millisecond 
    GtpRxMessageRate_o   => i_LRxGtpRxMessageRate,        -- : out std_logic_vector( 7 downto 0); -- Count per millisecond 

    -- Configuration signals
    -----------------------------
    --
    -- Source I/F configurations
    EnablePAER_i         => LRxPaerEn_i,                 -- in  std_logic;
    EnableHSSAER_i       => LRxHSSaerEn_i,               -- in  std_logic;
    EnableGTP_i          => LRxGtpEn_i,                  -- in  std_logic;
    EnableSPNNLNK_i      => LRxSpnnLnkEn_i,              -- in  std_logic;
    -- PAER
    RxPaerHighBits_i     => c_LRxPaerHighBits,           -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    PaerReqActLevel_i    => RxPaerReqActLevel_i,         -- in  std_logic;
    PaerAckActLevel_i    => RxPaerAckActLevel_i,         -- in  std_logic;
    PaerIgnoreFifoFull_i => RxPaerIgnoreFifoFull_i,      -- in  std_logic;
    PaerAckSetDelay_i    => RxPaerAckSetDelay_i,         -- in  std_logic_vector(7 downto 0);
    PaerSampleDelay_i    => RxPaerSampleDelay_i,         -- in  std_logic_vector(7 downto 0);
    PaerAckRelDelay_i    => RxPaerAckRelDelay_i,         -- in  std_logic_vector(7 downto 0);
    -- HSSAER
    RxSaerHighbits0_i    => c_LRxSaerHighBits0,          -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    RxSaerHighbits1_i    => c_LRxSaerHighBits1,          -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    RxSaerHighbits2_i    => c_LRxSaerHighBits2,          -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    RxSaerHighbits3_i    => c_LRxSaerHighBits3,          -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    HSSaerChanEn_i       => LRxSaerChanEn_i,             -- in  std_logic_vector(C_HSSAER_N_CHAN-1 downto 0);
    -- GTP
    RxGtpHighbits_i      => c_LRxGtpHighBits,            -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    -- SpiNNlink controls
    Spnn_start_key_i     => Spnn_start_key_i,            -- in  std_logic_vector(31 downto 0);
    Spnn_stop_key_i      => Spnn_stop_key_i,             -- in  std_logic_vector(31 downto 0);
    Spnn_cmd_start_o     => open,                        -- out std_logic;
    Spnn_cmd_stop_o      => open,                        -- out std_logic;
    Spnn_rx_mask_i       => Spnn_rx_mask_i,              -- in  std_logic_vector(31 downto 0);
    Spnn_keys_enable_i   => Spnn_ctrl_i(24),             -- in  std_logic;
    Spnn_parity_err_o    => Spnn_status_o(25),           -- out std_logic;
    Spnn_rx_err_o        => Spnn_status_o(24),           -- out std_logic; 
                        
    -- **********************************************
    -- Source Interfaces
    -- **********************************************

    -- Parallel AER
    -- ----------------------------------------------
    PAER_Addr_i          => i_LRxPaerAddr,               -- in  std_logic_vector(C_PAER_DSIZE-1 downto 0);
    PAER_Req_i           => i_LRxPaerReq,                -- in  std_logic;
    PAER_Ack_o           => i_LRxPaerAck,                -- out std_logic;

    -- HSSAER
    -- ----------------------------------------------
    HSSAER_Rx_i          => i_LRxHssaer,                -- in  std_logic_vector(0 to C_HSSAER_N_CHAN-1);

    -- GTP interface
    -- ----------------------------------------------
    RxGtpAlignRequest_o  => LRxRxGtpAlignRequest_o,            -- out std_logic;  
    
    -- GTP Wizard Interface
    -- Clock Ports
    GtpRxUsrClk2_i       => LRxGtpRxUsrClk2_i, 
    
    -- Reset FSM Control Ports
    SoftResetRx_o        => LRxSoftResetRx_o,                                
    GtpDataValid_o       => LRxGtpDataValid_o,                                
    
    -- -----------
    -- Receiver
    
    -- RX Initialization and Reset Ports
    GtpRxuserrdy_o       => LRxGtpRxuserrdy_o,                                      
    -- Receive Ports - FPGA RX Interface Ports 
    GtpRxdata_i          => LRxGtpRxdata_i,            
    -- Receive Ports - RX 8B/10B Decoder Ports 
    GtpRxchariscomma_i   => LRxGtpRxchariscomma_i,      
    GtpRxcharisk_i       => LRxGtpRxcharisk_i,          
    GtpRxdisperr_i       => LRxGtpRxdisperr_i,          
    GtpRxnotintable_i    => LRxGtpRxnotintable_i,       
    -- Receive Ports - RX Byte and Word Alignment Ports 
    GtpRxbyteisaligned_i => LRxGtpRxbyteisaligned_i,                           
    GtpRxbyterealign_i   => LRxGtpRxbyterealign_i,                            
    
    -- ------------ 
    -- Common ports
    GtpPllLock_i        => LRxGtpPllLock_i,                                        
    GtpPllRefclklost_i  => LRxGtpPllRefclklost_i,                                      

    -- SpiNNlink
    -- ----------------------------------------------
    data_2of7_from_spinnaker_i => i_LRxData2of7FromSpinnaker,
    ack_to_spinnaker_o         => i_LRxAckToSpinnaker,


    -- **********************************************
    -- Monitor interface
    -- **********************************************
    ToMonDataIn_o        => LRxData,               -- : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);  i_rxMonSrc(0).idx,      
    ToMonSrcRdy_o        => LRxSrcRdy,             -- : out std_logic;                                      i_rxMonSrc(0).vld,      
    ToMonDstRdy_i        => LRxDstRdy,             -- : in  std_logic;                                      i_rxMonDst(0).rdy,      
        
        
    -- **********************************************
    -- Debug signals
    -- **********************************************
    dbg_PaerDataOk       => open,                         -- out std_logic
    DBG_src_rdy          => open,
    DBG_dst_rdy          => open,
    DBG_err              => open, 
    DBG_run              => open,
    DBG_RX               => open,
    
    DBG_FIFO_0           => open,
    DBG_FIFO_1           => open,
    DBG_FIFO_2           => open,
    DBG_FIFO_3           => open,
    DBG_FIFO_4           => open                         
    );


u_rx_right_datapath : hpu_rx_datapath
  generic map (
    C_OUTPUT_DSIZE            => C_INTERNAL_DSIZE,
    C_PAER_DSIZE              => C_PAER_DSIZE,
    C_HAS_PAER                => C_RX_HAS_PAER,
    C_HAS_HSSAER              => C_RX_HAS_HSSAER,
    C_HSSAER_N_CHAN           => C_RX_HSSAER_N_CHAN,
    C_HAS_GTP                 => C_RX_HAS_GTP,
    C_GTP_DSIZE               => C_GTP_DSIZE,
    C_GTP_TXUSRCLK2_PERIOD_NS => C_GTP_TXUSRCLK2_PERIOD_NS,
    C_GTP_RXUSRCLK2_PERIOD_NS => C_GTP_RXUSRCLK2_PERIOD_NS,
    C_HAS_SPNNLNK             => C_RX_HAS_SPNNLNK,
    C_PSPNNLNK_WIDTH          => C_PSPNNLNK_WIDTH,
    C_SIM_TIME_COMPRESSION    => C_SIM_TIME_COMPRESSION
    )
  port map (

    -- **********************************************
    -- Barecontrol
    -- **********************************************
    -- Resets
    nRst                 => nRst,                        -- in  std_logic;
    -- System Clock domain
    Clk_i                => Clk_i,                    -- in  std_logic;
    En1Sec_i             => timing_i.en1s,-- : in  std_logic;
		-- HSSAER Clocks domain
		Clk_hs_p             => Clk_hs_p,                     -- in  std_logic;
		Clk_hs_n             => Clk_hs_n,                     -- in  std_logic;
    Clk_ls_p             => Clk_ls_p,                     -- in  std_logic;
    Clk_ls_n             => Clk_ls_n,                     -- in  std_logic;
 
 
    -- **********************************************
    -- Controls
    -- **********************************************
    --
    -- In case of aux channel the HPU header is 
    -- adapted to what received
    -- ----------------------------------------------
    Aux_Channel_i        => '0',


    -- **********************************************
    -- uController Interface
    -- **********************************************

    -- Control signals
    -- ----------------------------------------------
    PaerFlushFifos_i     => RRxPaerFlushFifos_i,         -- in  std_logic;
    
    -- Status signals
    -----------------------------
    PaerFifoFull_o       => RRxPaerFifoFull_o,           -- out std_logic;
    RxSaerStat_o         => RRxSaerStat_o,               -- out t_RxSaerStat_array(C_HSSAER_N_CHAN-1 downto 0);
    RxGtpStat_o          => RRxGtpStat_o,                -- out t_RxGtpStat;
    RxSpnnlnkStat_o      => RRxSpnnlnkStat_o,            -- out t_RxSpnnlnkStat;
    
    -- GTP Statistics        
    GtpRxDataRate_o      => i_RRxGtpRxDataRate,          -- : out std_logic_vector(15 downto 0); -- Count per millisecond 
    GtpRxAlignRate_o     => i_RRxGtpRxAlignRate,         -- : out std_logic_vector( 7 downto 0); -- Count per millisecond 
    GtpRxMsgRate_o       => i_RRxGtpRxMsgRate,           -- : out std_logic_vector(15 downto 0); -- Count per millisecond 
    GtpRxIdleRate_o      => i_RRxGtpRxIdleRate,          -- : out std_logic_vector(15 downto 0); -- Count per millisecond 
    GtpRxEventRate_o     => i_RRxGtpRxEventRate,         -- : out std_logic_vector(15 downto 0); -- Count per millisecond 
    GtpRxMessageRate_o   => i_RRxGtpRxMessageRate,       -- : out std_logic_vector( 7 downto 0); -- Count per millisecond 

    -- Configuration signals
    -----------------------------
    --
    -- Source I/F configurations
    EnablePAER_i         => RRxPaerEn_i,                 -- in  std_logic;
    EnableHSSAER_i       => RRxHSSaerEn_i,               -- in  std_logic;
    EnableGTP_i          => RRxGtpEn_I,                  -- in  std_logic;
    EnableSPNNLNK_i      => RRxSpnnLnkEn_i,              -- in  std_logic;
    -- PAER
    RxPaerHighBits_i     => c_RRxPaerHighBits,           -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    PaerReqActLevel_i    => RxPaerReqActLevel_i,         -- in  std_logic;
    PaerAckActLevel_i    => RxPaerAckActLevel_i,         -- in  std_logic;
    PaerIgnoreFifoFull_i => RxPaerIgnoreFifoFull_i,      -- in  std_logic;
    PaerAckSetDelay_i    => RxPaerAckSetDelay_i,         -- in  std_logic_vector(7 downto 0);
    PaerSampleDelay_i    => RxPaerSampleDelay_i,         -- in  std_logic_vector(7 downto 0);
    PaerAckRelDelay_i    => RxPaerAckRelDelay_i,         -- in  std_logic_vector(7 downto 0);
    -- HSSAER
    RxSaerHighbits0_i    => c_RRxSaerHighBits0,          -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    RxSaerHighbits1_i    => c_RRxSaerHighBits1,          -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    RxSaerHighbits2_i    => c_RRxSaerHighBits2,          -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    RxSaerHighbits3_i    => c_RRxSaerHighBits3,          -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    HSSaerChanEn_i       => RRxSaerChanEn_i,             -- in  std_logic_vector(C_HSSAER_N_CHAN-1 downto 0);
    -- GTP
    RxGtpHighbits_i      => c_RRxGtpHighBits,            -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    -- SpiNNlink controls
    Spnn_start_key_i     => Spnn_start_key_i,            -- in  std_logic_vector(31 downto 0);
    Spnn_stop_key_i      => Spnn_stop_key_i,             -- in  std_logic_vector(31 downto 0);
    Spnn_cmd_start_o     => open,                        -- out std_logic;
    Spnn_cmd_stop_o      => open,                        -- out std_logic;
    Spnn_rx_mask_i       => Spnn_rx_mask_i,              -- in  std_logic_vector(31 downto 0);
    Spnn_keys_enable_i   => Spnn_ctrl_i(16),             -- in  std_logic;
    Spnn_parity_err_o    => Spnn_status_o(17),           -- out std_logic;
    Spnn_rx_err_o        => Spnn_status_o(16),           -- out std_logic;
                        
    -- **********************************************
    -- Source Interfaces
    -- **********************************************

    -- Parallel AER
    -- ----------------------------------------------
    PAER_Addr_i          => i_RRxPaerAddr,             -- in  std_logic_vector(C_PAER_DSIZE-1 downto 0);
    PAER_Req_i           => i_RRxPaerReq,              -- in  std_logic;
    PAER_Ack_o           => i_RRxPaerAck,              -- out std_logic;

    -- HSSAER
    -- ----------------------------------------------
    HSSAER_Rx_i          => i_RRxHssaer,                -- in  std_logic_vector(0 to C_HSSAER_N_CHAN-1);

    -- GTP interface
    -- ----------------------------------------------
    RxGtpAlignRequest_o  => RRxRxGtpAlignRequest_o,            -- out std_logic;  
    
    -- GTP Wizard Interface
    -- Clock Ports
    GtpRxUsrClk2_i       => RRxGtpRxUsrClk2_i, 
    
    -- Reset FSM Control Ports
    SoftResetRx_o        => RRxSoftResetRx_o,                                
    GtpDataValid_o       => RRxGtpDataValid_o,                                

    -- -----------
    -- Receiver
    
    -- RX Initialization and Reset Ports
    GtpRxuserrdy_o       => RRxGtpRxuserrdy_o,                                           
    -- Receive Ports - FPGA RX Interface Ports 
    GtpRxdata_i          => RRxGtpRxdata_i,            
    -- Receive Ports - RX 8B/10B Decoder Ports 
    GtpRxchariscomma_i   => RRxGtpRxchariscomma_i,      
    GtpRxcharisk_i       => RRxGtpRxcharisk_i,          
    GtpRxdisperr_i       => RRxGtpRxdisperr_i,          
    GtpRxnotintable_i    => RRxGtpRxnotintable_i,       
    -- Receive Ports - RX Byte and Word Alignment Ports 
    GtpRxbyteisaligned_i => RRxGtpRxbyteisaligned_i,                           
    GtpRxbyterealign_i   => RRxGtpRxbyterealign_i,                            
    
    -- ------------ 
    -- Common ports
    GtpPllLock_i         => RRxGtpPllLock_i,                                        
    GtpPllRefclklost_i   => RRxGtpPllRefclklost_i,                                      

    -- SpiNNlink
    -- ----------------------------------------------
    data_2of7_from_spinnaker_i => i_RRxData2of7FromSpinnaker,
    ack_to_spinnaker_o         => i_RRxAckToSpinnaker,


    -- **********************************************
    -- Monitor interface
    -- **********************************************
    ToMonDataIn_o        => RRxData,               -- : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);  i_rxMonSrc(1).idx,      
    ToMonSrcRdy_o        => RRxSrcRdy,             -- : out std_logic;                                      i_rxMonSrc(1).vld,      
    ToMonDstRdy_i        => RRxDstRdy,             -- : in  std_logic;                                      i_rxMonDst(1).rdy,      
        
        
    -- **********************************************
    -- Debug signals
    -- **********************************************
    dbg_PaerDataOk       => open,                         -- out std_logic
    DBG_src_rdy          => open,
    DBG_dst_rdy          => open,
    DBG_err              => open, 
    DBG_run              => open,
    DBG_RX               => open,
    
    DBG_FIFO_0           => open,
    DBG_FIFO_1           => open,
    DBG_FIFO_2           => open,
    DBG_FIFO_3           => open,
    DBG_FIFO_4           => open                         
    );


u_rx_aux_datapath : hpu_rx_datapath
  generic map (
    C_OUTPUT_DSIZE            => C_INTERNAL_DSIZE,
    C_PAER_DSIZE              => C_PAER_DSIZE,
    C_HAS_PAER                => C_RX_HAS_PAER,
    C_HAS_HSSAER              => C_RX_HAS_HSSAER,
    C_HSSAER_N_CHAN           => C_RX_HSSAER_N_CHAN,
    C_HAS_GTP                 => C_RX_HAS_GTP,
    C_GTP_DSIZE               => C_GTP_DSIZE,
    C_GTP_TXUSRCLK2_PERIOD_NS => C_GTP_TXUSRCLK2_PERIOD_NS,
    C_GTP_RXUSRCLK2_PERIOD_NS => C_GTP_RXUSRCLK2_PERIOD_NS,
    C_HAS_SPNNLNK             => C_RX_HAS_SPNNLNK,
    C_PSPNNLNK_WIDTH          => C_PSPNNLNK_WIDTH,
    C_SIM_TIME_COMPRESSION    => C_SIM_TIME_COMPRESSION
    )
  port map (

    -- **********************************************
    -- Barecontrol
    -- **********************************************
    -- Resets
    nRst                 => nRst,                         -- in  std_logic;
    -- System Clock domain
    Clk_i                => Clk_i,                        -- in  std_logic;
    En1Sec_i             => timing_i.en1s,                -- : in  std_logic;
		-- HSSAER Clocks domain
		Clk_hs_p             => Clk_hs_p,                     -- in  std_logic;
		Clk_hs_n             => Clk_hs_n,                     -- in  std_logic;
    Clk_ls_p             => Clk_ls_p,                     -- in  std_logic;
    Clk_ls_n             => Clk_ls_n,                     -- in  std_logic;
 
 
    -- **********************************************
    -- Controls
    -- **********************************************
    --
    -- In case of aux channel the HPU header is 
    -- adapted to what received
    -- ----------------------------------------------
    Aux_Channel_i        => '1',


    -- **********************************************
    -- uController Interface
    -- **********************************************

    -- Control signals
    -- ----------------------------------------------
    PaerFlushFifos_i     => AuxRxPaerFlushFifos_i,         -- in  std_logic;
    
    -- Status signals
    -----------------------------
    PaerFifoFull_o       => AuxRxPaerFifoFull_o,           -- out std_logic;
    RxSaerStat_o         => AuxRxSaerStat_o,               -- out t_RxSaerStat_array(C_HSSAER_N_CHAN-1 downto 0);
    RxGtpStat_o          => AuxRxGtpStat_o,                -- out t_RxGtpStat;
    RxSpnnlnkStat_o      => AuxRxSpnnlnkStat_o,            -- out t_RxSpnnlnkStat;
    
    -- GTP Statistics        
    GtpRxDataRate_o      => i_AuxRxGtpRxDataRate,          -- : out std_logic_vector(15 downto 0); -- Count per millisecond 
    GtpRxAlignRate_o     => i_AuxRxGtpRxAlignRate,         -- : out std_logic_vector( 7 downto 0); -- Count per millisecond 
    GtpRxMsgRate_o       => i_AuxRxGtpRxMsgRate,           -- : out std_logic_vector(15 downto 0); -- Count per millisecond 
    GtpRxIdleRate_o      => i_AuxRxGtpRxIdleRate,          -- : out std_logic_vector(15 downto 0); -- Count per millisecond 
    GtpRxEventRate_o     => i_AuxRxGtpRxEventRate,         -- : out std_logic_vector(15 downto 0); -- Count per millisecond 
    GtpRxMessageRate_o   => i_AuxRxGtpRxMessageRate,       -- : out std_logic_vector( 7 downto 0); -- Count per millisecond 

    -- Configuration signals
    -----------------------------
    --
    -- Source I/F configurations
    EnablePAER_i         => AuxRxPaerEn_i,                 -- in  std_logic;
    EnableHSSAER_i       => AuxRxHSSaerEn_i,               -- in  std_logic;
    EnableGTP_i          => AuxRxGtpEn_I,                  -- in  std_logic;
    EnableSPNNLNK_i      => AuxRxSpnnLnkEn_i,              -- in  std_logic;
    -- PAER
    RxPaerHighBits_i     => c_AuxRxPaerHighBits,           -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    PaerReqActLevel_i    => RxPaerReqActLevel_i,         -- in  std_logic;
    PaerAckActLevel_i    => RxPaerAckActLevel_i,         -- in  std_logic;
    PaerIgnoreFifoFull_i => RxPaerIgnoreFifoFull_i,      -- in  std_logic;
    PaerAckSetDelay_i    => RxPaerAckSetDelay_i,         -- in  std_logic_vector(7 downto 0);
    PaerSampleDelay_i    => RxPaerSampleDelay_i,         -- in  std_logic_vector(7 downto 0);
    PaerAckRelDelay_i    => RxPaerAckRelDelay_i,         -- in  std_logic_vector(7 downto 0);
    -- HSSAER
    RxSaerHighbits0_i    => c_AuxRxSaerHighBits0,          -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    RxSaerHighbits1_i    => c_AuxRxSaerHighBits1,          -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    RxSaerHighbits2_i    => c_AuxRxSaerHighBits2,          -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    RxSaerHighbits3_i    => c_AuxRxSaerHighBits3,          -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    HSSaerChanEn_i       => AuxRxSaerChanEn_i,             -- in  std_logic_vector(C_HSSAER_N_CHAN-1 downto 0);
    -- GTP
    RxGtpHighbits_i      => c_AuxRxGtpHighBits,            -- in  std_logic_vector(C_INTERNAL_DSIZE-1 downto C_PAER_DSIZE);
    -- SpiNNlink controls
    Spnn_start_key_i     => Spnn_start_key_i,            -- in  std_logic_vector(31 downto 0);
    Spnn_stop_key_i      => Spnn_stop_key_i,             -- in  std_logic_vector(31 downto 0);
    Spnn_cmd_start_o     => open,                        -- out std_logic;
    Spnn_cmd_stop_o      => open,                        -- out std_logic;
    Spnn_rx_mask_i       => Spnn_rx_mask_i,              -- in  std_logic_vector(31 downto 0);
    Spnn_keys_enable_i   => Spnn_ctrl_i(8),             -- in  std_logic;
    Spnn_parity_err_o    => Spnn_status_o(9),           -- out std_logic;
    Spnn_rx_err_o        => Spnn_status_o(8),           -- out std_logic;
                        
    -- **********************************************
    -- Source Interfaces
    -- **********************************************

    -- Parallel AER
    -- ----------------------------------------------
    PAER_Addr_i          => i_AuxRxPaerAddr,             -- in  std_logic_vector(C_PAER_DSIZE-1 downto 0);
    PAER_Req_i           => i_AuxRxPaerReq,              -- in  std_logic;
    PAER_Ack_o           => i_AuxRxPaerAck,              -- out std_logic;

    -- HSSAER
    -- ----------------------------------------------
    HSSAER_Rx_i          => i_AuxRxHssaer,                -- in  std_logic_vector(0 to C_HSSAER_N_CHAN-1);

    -- GTP interface
    -- ----------------------------------------------
    RxGtpAlignRequest_o  => AuxRxRxGtpAlignRequest_o,            -- out std_logic;  
    
    -- GTP Wizard Interface
    -- Clock Ports
    GtpRxUsrClk2_i       => AuxRxGtpRxUsrClk2_i, 
    
    -- Reset FSM Control Ports
    SoftResetRx_o        => AuxRxSoftResetRx_o,                                
    GtpDataValid_o       => AuxRxGtpDataValid_o,                                
    
    -- -----------
    -- Receiver
    
    -- RX Initialization and Reset Ports
    GtpRxuserrdy_o       => AuxRxGtpRxuserrdy_o,                                           
    -- Receive Ports - FPGA RX Interface Ports 
    GtpRxdata_i          => AuxRxGtpRxdata_i,            
    -- Receive Ports - RX 8B/10B Decoder Ports 
    GtpRxchariscomma_i   => AuxRxGtpRxchariscomma_i,      
    GtpRxcharisk_i       => AuxRxGtpRxcharisk_i,          
    GtpRxdisperr_i       => AuxRxGtpRxdisperr_i,          
    GtpRxnotintable_i    => AuxRxGtpRxnotintable_i,       
    -- Receive Ports - RX Byte and Word Alignment Ports 
    GtpRxbyteisaligned_i => AuxRxGtpRxbyteisaligned_i,                           
    GtpRxbyterealign_i   => AuxRxGtpRxbyterealign_i,                            
    
    -- ------------ 
    -- Common ports
    GtpPllLock_i        => AuxRxGtpPllLock_i,                                        
    GtpPllRefclklost_i  => AuxRxGtpPllRefclklost_i,                                      

    -- SpiNNlink
    -- ----------------------------------------------
    data_2of7_from_spinnaker_i => i_AuxRxData2of7FromSpinnaker,
    ack_to_spinnaker_o         => i_AuxRxAckToSpinnaker,


    -- **********************************************
    -- Monitor interface
    -- **********************************************
    ToMonDataIn_o        => AuxRxData,               -- : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);  i_rxMonSrc(2).idx,      
    ToMonSrcRdy_o        => AuxRxSrcRdy,             -- : out std_logic;                                      i_rxMonSrc(2).vld,      
    ToMonDstRdy_i        => AuxRxDstRdy,             -- : in  std_logic;                                      i_rxMonDst(2).rdy,      
        
        
    -- **********************************************
    -- Debug signals
    -- **********************************************
    dbg_PaerDataOk       => open,                         -- out std_logic
    DBG_src_rdy          => open,
    DBG_dst_rdy          => open,
    DBG_err              => open, 
    DBG_run              => open,
    DBG_RX               => open,
    
    DBG_FIFO_0           => open,
    DBG_FIFO_1           => open,
    DBG_FIFO_2           => open,
    DBG_FIFO_3           => open,
    DBG_FIFO_4           => open                         
    );



--Interceptions
---------------------

LEFT_INTERCEPTION_TRUE_gen: if C_RX_LEFT_INTERCEPTION = true generate
begin
    LRxData_o           <= LRxData;
    LRxSrcRdy_o         <= LRxSrcRdy;
    LRxDstRdy           <= LRxDstRdy_i;
    i_rxMonSrc(0).idx   <= LRxBypassData_i;
    i_rxMonSrc(0).vld   <= LRxBypassSrcRdy_i; 
    LRxBypassDstRdy_o   <= i_rxMonDst(0).rdy;
end generate;
LEFT_INTERCEPTION_FALSE_gen: if C_RX_LEFT_INTERCEPTION = false generate
begin
    i_rxMonSrc(0).idx   <= LRxData;
    i_rxMonSrc(0).vld   <= LRxSrcRdy; 
    LRxDstRdy           <= i_rxMonDst(0).rdy;
end generate;


RIGHT_INTERCEPTION_TRUE_gen: if C_RX_RIGHT_INTERCEPTION = true generate
begin
    RRxData_o           <= RRxData;
    RRxSrcRdy_o         <= RRxSrcRdy;
    RRxDstRdy           <= RRxDstRdy_i;
    i_rxMonSrc(1).idx   <= RRxBypassData_i;
    i_rxMonSrc(1).vld   <= RRxBypassSrcRdy_i; 
    RRxBypassDstRdy_o   <= i_rxMonDst(1).rdy;  
end generate;
RIGHT_INTERCEPTION_FALSE_gen: if C_RX_RIGHT_INTERCEPTION = false generate
begin
    i_rxMonSrc(1).idx   <= RRxData;
    i_rxMonSrc(1).vld   <= RRxSrcRdy; 
    RRxDstRdy           <= i_rxMonDst(1).rdy;
end generate;


AUX_INTERCEPTION_TRUE_gen: if C_RX_AUX_INTERCEPTION = true generate
begin
    AuxRxData_o         <= AuxRxData;
    AuxRxSrcRdy_o       <= AuxRxSrcRdy;
    AuxRxDstRdy         <= AuxRxDstRdy_i;
    i_rxMonSrc(2).idx   <= AuxRxBypassData_i;
    i_rxMonSrc(2).vld   <= AuxRxBypassSrcRdy_i; 
    AuxRxBypassDstRdy_o <= i_rxMonDst(2).rdy;  
end generate;
AUX_INTERCEPTION_FALSE_gen: if C_RX_AUX_INTERCEPTION = false generate
begin
    i_rxMonSrc(2).idx   <= AuxRxData;
    i_rxMonSrc(2).vld   <= AuxRxSrcRdy; 
    AuxRxDstRdy         <= i_rxMonDst(2).rdy;
end generate;

--        ToMonDataIn_o        => RRxData_o,               -- : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);  i_rxMonSrc(1).idx, 
--        ToMonSrcRdy_o        => RRxSrcRdy_o,             -- : out std_logic;                                      i_rxMonSrc(1).vld, 
--        ToMonDstRdy_i        => RRxDstRdy_i,             -- : in  std_logic;                                      i_rxMonDst(1).rdy, 
       
--        RRxData_o               : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
--        RRxSrcRdy_o             : out std_logic;
--        RRxDstRdy_i             : in  std_logic;
--        RRxBypassData_i         : in  std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
--        RRxBypassSrcRdy_i       : in  std_logic;
--        RRxBypassDstRdy_o       : out std_logic;
--        --
--        LRxData_o               : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
--        LRxSrcRdy_o             : out std_logic;
--        LRxDstRdy_i             : in  std_logic;
--        LRxBypassData_i         : in  std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
--        LRxBypassSrcRdy_i       : in  std_logic;
--        LRxBypassDstRdy_o       : out std_logic;
--        --
--        AuxRxData_o             : out std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
--        AuxRxSrcRdy_o           : out std_logic;
--        AuxRxDstRdy_i           : in  std_logic;
--        AuxRxBypassData_i       : in  std_logic_vector(C_INTERNAL_DSIZE-1 downto 0);
--        AuxRxBypassSrcRdy_i     : in  std_logic;
--        AuxRxBypassDstRdy_o     : out std_logic;            
        

    u_RxArbiter : neuserial_PAER_arbiter
        generic map (
            C_NUM_CHAN     => 3,
            C_ODATA_WIDTH  => 32
        )
        port map (
            Clk                => Clk_i,                  -- in  std_logic;
            nRst               => nRst,                      -- in  std_logic;

            SplittedPaerSrc_i  => i_rxMonSrc,                -- in  t_PaerSrc_array(0 to C_NUM_CHAN-1);
            SplittedPaerDst_o  => i_rxMonDst,                -- out t_PaerDst_array(0 to C_NUM_CHAN-1);

            PaerData_o         => i_rxMonData,               -- out std_logic_vector(31 downto 0);
            PaerSrcRdy_o       => i_rxMonSrcRdy,             -- out std_logic;
            PaerDstRdy_i       => i_rxMonDstRdy              -- in  std_logic
        );


   
    ---------------------
    -- Loopbacks
    ---------------------

    -- Local Near and Remote Loopback

    i_monData   <= i_seqData   when LocNearLoopback_i = '1' else
                   i_rxMonData;
    i_monSrcRdy <= i_seqSrcRdy when LocNearLoopback_i = '1' else
                   i_rxMonSrcRdy;

    i_seqDstRdy <= i_monDstRdy when LocNearLoopback_i = '1' else
                   '1'         when RemoteLoopback_i  = '1' else
                   i_txSeqDstRdy;

    i_rxMonDstRdy <= i_txSeqDstRdy when RemoteLoopback_i  = '1' else
                     '1'           when LocNearLoopback_i = '1' else
                     i_monDstRdy;

    i_txSeqData   <= i_rxMonData   when RemoteLoopback_i = '1' else
                     i_seqData;
    i_txSeqSrcRdy <= i_rxMonSrcRdy when RemoteLoopback_i = '1' else
                     i_seqSrcRdy;


    -------------------------------
    -- Sequencer & Monitor core
    -------------------------------

    u_CoreMonSeqRR : CoreMonSeqRR
        generic map (
            C_PAER_DSIZE                         => C_PAER_DSIZE,
            TestEnableSequencerNoWait            => c_TestEnableSequencerNoWait,
            TestEnableSequencerToMonitorLoopback => c_TestEnableSequencerToMonitorLoopback,
            EnableMonitorControlsSequencerToo    => c_EnableMonitorControlsSequencerToo
        )
        port map (
            Reset_xRBI              => nRst,                     -- in  std_logic;
            CoreClk_xCI             => Clk_i,                 -- in  std_logic;
            --
            FlushRXFifos_xSI        => FlushRXFifos_i,           -- in  std_logic;
            FlushTXFifos_xSI        => FlushTXFifos_i,           -- in  std_logic;
            --ChipType_xSI            => ChipType,                 -- in  std_logic;
            DmaLength_xDI           => DmaLength_i,              -- in  std_logic_vector(15 downto 0);
            --
            Timing_xSI              => timing_i,                 -- in  time_tick;
            --
            MonInAddr_xDI           => i_monData,                -- in  std_logic_vector(31 downto 0);
            MonInSrcRdy_xSI         => i_monSrcRdy,              -- in  std_logic;
            MonInDstRdy_xSO         => i_monDstRdy,              -- out std_logic;
            --
            SeqOutAddr_xDO          => i_seqData,                -- out std_logic_vector(31 downto 0);
            SeqOutSrcRdy_xSO        => i_seqSrcRdy,              -- out std_logic;
            SeqOutDstRdy_xSI        => i_seqDstRdy,              -- in  std_logic;
            -- Time stamper
            CleanTimer_xSI          => CleanTimer_i,             -- in  std_logic;
            WrapDetected_xSO        => WrapDetected_o,           -- out std_logic;
            FullTimestamp_i         => FullTimestamp_i,          -- in  std_logic;  
            --
            EnableMonitor_xSI       => '1',                      -- in  std_logic;
            CoreReady_xSI           => '1',                      -- in  std_logic;
            --
            TxTSMode_xDI            => TxTSMode_i,               -- in  std_logic_vector(1 downto 0);
            TxTSTimeoutSel_xDI      => TxTSTimeoutSel_i,         -- in  std_logic_vector(3 downto 0);
            TxTSRetrigCmd_xSI       => TxTSRetrigCmd_i,          -- in  std_logic;
            TxTSRearmCmd_xSI        => TxTSRearmCmd_i,           -- in  std_logic;
            TxTSRetrigStatus_xSO    => TxTSRetrigStatus_o,       -- out std_logic;
            TxTSTimeoutCounts_xSO   => TxTSTimeoutCounts_o,      -- out std_logic;
            TxTSMaskSel_xSI         => TxTSMaskSel_i,            -- in  std_logic_vector(1 downto 0);
            --
            FifoCoreDat_xDO         => FifoCoreDat_o,            -- out std_logic_vector(31 downto 0);
            FifoCoreRead_xSI        => FifoCoreRead_i,           -- in  std_logic;
            FifoCoreEmpty_xSO       => FifoCoreEmpty_o,          -- out std_logic;
            FifoCoreAlmostEmpty_xSO => FifoCoreAlmostEmpty_o,    -- out std_logic;
            FifoCoreBurstReady_xSO  => FifoCoreBurstReady_o,     -- out std_logic;
            FifoCoreFull_xSO        => FifoCoreFull_o,           -- out std_logic;
            FifoCoreNumData_o       => FifoCoreNumData_o,        -- out std_logic_vector(10 downto 0);
            --
            CoreFifoDat_xDI         => CoreFifoDat_i,            -- in  std_logic_vector(31 downto 0);
            CoreFifoWrite_xSI       => CoreFifoWrite_i,          -- in  std_logic;
            CoreFifoFull_xSO        => CoreFifoFull_o,           -- out std_logic;
            CoreFifoAlmostFull_xSO  => CoreFifoAlmostFull_o,     -- out std_logic;
            CoreFifoEmpty_xSO       => CoreFifoEmpty_o,          -- out std_logic;
            --
            --BiasFinished_xSO        => BiasFinished,             -- out std_logic;
            --ClockLow_xDI            => ClockLow,                 -- in  natural;
            --LatchTime_xDI           => LatchTime,                -- in  natural;
            --SetupHold_xDI           => SetupHold,                -- in  natural;
            --PrescalerValue_xDI      => PrescalerValue,           -- in  std_logic_vector(31 downto 0);
            --BiasProgPins_xDO        => i_BiasProgPins_xD,        -- out std_logic_vector(7 downto 0);
            ---------------------------------------------------------------------------
            -- Output neurons threshold
            --OutThresholdVal_xDI     => OutThresholdVal           -- in  std_logic_vector(31 downto 0)
            DBG_din             => DBG_din,   
            DBG_wr_en           => DBG_wr_en,       
            DBG_rd_en           => DBG_rd_en,       
            DBG_dout            => DBG_dout,            
            DBG_full            => DBG_full,        
            DBG_almost_full     => DBG_almost_full, 
            DBG_overflow        => DBG_overflow,      
            DBG_empty           => DBG_empty,            
            DBG_almost_empty    => DBG_almost_empty,
            DBG_underflow       => DBG_underflow,   
            DBG_data_count      => DBG_data_count,
            DBG_Timestamp_xD    => DBG_Timestamp_xD,
            DBG_MonInAddr_xD    => DBG_MonInAddr_xD, 
            DBG_MonInSrcRdy_xS  => DBG_MonInSrcRdy_xS,
            DBG_MonInDstRdy_xS  => DBG_MonInDstRdy_xS,
            DBG_RESETFIFO       => DBG_RESETFIFO
 
 
        );




    -----------------------------------------------------------------------------
    -- LEDs
    -----------------------------------------------------------------------------
    LEDo_o <= '1';
    LEDr_o <= '1';
    LEDy_o <= '1';
    
    DBG_CH0_DATA <= i_rxMonSrc(0).idx;
    DBG_CH0_SRDY <= i_rxMonSrc(0).vld;
    DBG_CH0_DRDY <= i_rxMonDst(0).rdy;

    DBG_CH1_DATA <= i_rxMonSrc(1).idx;
    DBG_CH1_SRDY <= i_rxMonSrc(1).vld;
    DBG_CH1_DRDY <= i_rxMonDst(1).rdy;

    DBG_CH2_DATA <= i_rxMonSrc(2).idx;
    DBG_CH2_SRDY <= i_rxMonSrc(2).vld;
    DBG_CH2_DRDY <= i_rxMonDst(2).rdy;
    


end architecture str;

-------------------------------------------------------------------------------
