library ieee;
    use ieee.std_logic_1164.all;
    use ieee.numeric_std.all;

library datapath;
    use datapath.constants.all;
    use datapath.types.all;
    
library swissknife;
    use swissknife.types.all;

package components is
 
end package components;
